`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/11/09 20:35:47
// Design Name: 
// Module Name: tb_cpu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_cpu();
reg         clk,rst,en_in,en_ram_out;
reg  [15:0] ins;
wire        en_ram_in;
wire [15:0] addr;

cpu test_cpu(
    .clk (clk),
    .rst (rst),
    .en_in (en_in),
    .en_ram_in (en_ram_in), 
    .ins (ins),	
    .en_ram_out (en_ram_out),
    .addr (addr)   	
);

parameter Tclk = 10;

initial begin
	    //define clk
	    clk = 0;
        forever #(Tclk/2) clk = ~clk;
		end
        
initial begin
		//define rst
		rst = 0;
		#(Tclk*4) rst = 1;
		end

initial begin                
		//define en_in and en_ram_out
		en_in = 0;
		en_ram_out = 0;
		#(Tclk*8) en_in = 1;//enabling state_transition
		#(Tclk*2) en_ram_out = 1;//anabling ir
end

initial begin
         //define ins ,you can assign 0000_0000_0000_0001
		    //0000_0100_0000_0010 and so on to ins.
		           ins = 16'b0000_0000_0000_0000;

	    #(Tclk*10)  ins = 16'b0011_0000_0000_0000; //MOV（0000000000001000）
	    #(Tclk*10)  ins = 16'b0011_0000_1000_0100; //MOV (0000000000000100(im))
	    
	    #(Tclk*10)  ins = 16'b1100_0001_0000_0000; //ls（0000000000010000）
	    
        #(Tclk*10)  ins = 16'b1101_0001_0000_0000; //rs (0000000000010000)
        
        #(Tclk*10)  ins = 16'b1001_0000_0000_0000; //AND（1111111111111111&0000000000001000）
        #(Tclk*10)  ins = 16'b1001_0000_1000_0100; //AND (1111111111111111&0000000000000100(im))
            
        #(Tclk*10)  ins = 16'b1010_0000_0000_0000; //OR（1111111111111111|0000000000001000）
        #(Tclk*10)  ins = 16'b1010_0000_1000_0100; //OR (1111111111111111|0000000000000100(im))
        
	    #(Tclk*10)  ins = 16'b0100_0000_0000_0000; //ADD（1111111111111111+0000000000001000,carryout）
	    #(Tclk*10)  ins = 16'b0100_0000_1000_0100; //ADD (1111111111111111+0000000000000100(im),carryout)
	    #(Tclk*10)  ins = 16'b0100_0001_0000_0000; //ADD（000000000010000+0000000010000000）
        #(Tclk*10)  ins = 16'b0100_0001_1000_0100; //ADD (000000000010000+0000000000000100(im))
        
        #(Tclk*10)  ins = 16'b0101_0000_0000_0000; //SUB（1111111111111111-0000000000001000）
        #(Tclk*10)  ins = 16'b0101_0000_1000_0100; //SUB (1111111111111111-0000000000000100(im))
        #(Tclk*10)  ins = 16'b0101_0001_0000_0000; //SUB（000000000010000-0000000010000000,carryout）
        #(Tclk*10)  ins = 16'b0101_0001_1010_0000; //SUB (000000000010000-0000000000100000(im),carryout)
        
	    #(Tclk*10)  ins = 16'b1011_0000_0000_0000; //compare(1111111111111111>0000000000001000)
	    #(Tclk*10)  ins = 16'b1011_0000_1000_1001; //compare(1111111111111111>0000000000001001(im))
	    #(Tclk*10)  ins = 16'b1011_0001_0000_0000; //compare（000000000010000<0000000010000000）
        #(Tclk*10)  ins = 16'b1011_0001_1010_0000; //compare (000000000010000<0000000000100000(im))
	  	#(Tclk*10)  ins = 16'b1011_0010_0000_0000; //compare（000000000000100=0000000000000100）
        #(Tclk*10)  ins = 16'b1011_0010_1000_0100; //compare (000000000000100=0000000000000100(im))
        
        #(Tclk*10)  ins = 16'b0110_0000_0000_0000; //MUL（1111111111111111*0000000000001000,carryout）
        #(Tclk*10)  ins = 16'b0110_0000_1000_0100; //MUL (1111111111111111*0000000000000100(im),carryout)     
        #(Tclk*10)  ins = 16'b0110_0001_0000_0000; //MUL（000000000010000*0000000010000000）
        #(Tclk*10)  ins = 16'b0110_0001_1000_0100; //MUL (000000000010000*0000000000000100(im))
       
        #(Tclk*10)  ins = 16'b0111_0000_0000_0000; //DIV（1111111111111111/0000000000001000）
        #(Tclk*10)  ins = 16'b0111_0000_1000_0100; //DIV (1111111111111111/0000000000000100(im))
        #(Tclk*10)  ins = 16'b0111_0001_0000_0000; //DIV（000000000010000/0000000010000000）
        #(Tclk*10)  ins = 16'b0111_0001_1010_0000; //DIV (000000000010000/0000000000100000(im))
       
       	#(Tclk*10)  ins = 16'b1100_0001_0000_0000; //ls（0000000000010000）
       	
     // #(Tclk*10)  ins = 16'b1110_0001_0000_0000; //rs (0000000000010000)
       	
	    #(Tclk*6)  en_in = 0;  en_ram_out = 0;
	    
        end
       
initial begin
    #(Tclk*400)  $stop;
end

endmodule
